* Classical
.include TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param length=2u

.param width_12={40u}
.param width_34={30u}
.param width_58={9u}
.param width_6={200u}
.param width_7={28u}

.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
Iref gnd ref 24u
vinp inp gnd dc 0.9 ac 0.05m sin(0.9 0.05m 10k 0 0 0) 
vinn inn gnd dc 0.9 ac -0.05m sin(0.9 -0.05m 10k 0 0 0)

CL out gnd 1p
Cc k out 1p
Rz d2 k 2.2k

M1      d1     inn      d5     gnd  CMOSN   W={width_12}   L={2*length}
+ AS={5*width_12*LAMBDA} PS={10*LAMBDA+2*width_12} AD={5*width_12*LAMBDA} PD={10*LAMBDA+2*width_12}
M2      d2     inp      d5     gnd  CMOSN   W={width_12}   L={2*length}
+ AS={5*width_12*LAMBDA} PS={10*LAMBDA+2*width_12} AD={5*width_12*LAMBDA} PD={10*LAMBDA+2*width_12}
M3      d1     d1       vdd    vdd  CMOSP   W={width_34}   L={length}
+ AS={5*width_34*LAMBDA} PS={10*LAMBDA+2*width_34} AD={5*width_34*LAMBDA} PD={10*LAMBDA+2*width_34}
M4      d2     d1       vdd    vdd  CMOSP   W={width_34}   L={length}
+ AS={5*width_34*LAMBDA} PS={10*LAMBDA+2*width_34} AD={5*width_34*LAMBDA} PD={10*LAMBDA+2*width_34}
M5      d5     ref      gnd    gnd  CMOSN   W={width_58}   L={length}
+ AS={5*width_58*LAMBDA} PS={10*LAMBDA+2*width_58} AD={5*width_58*LAMBDA} PD={10*LAMBDA+2*width_58}
M6      out    d2       vdd    vdd  CMOSP   W={width_6}   L={length}
+ AS={5*width_6*LAMBDA} PS={10*LAMBDA+2*width_6} AD={5*width_6*LAMBDA} PD={10*LAMBDA+2*width_6}
M7      out    ref      gnd     gnd  CMOSN   W={width_7}   L={length}
+ AS={5*width_7*LAMBDA} PS={10*LAMBDA+2*width_7} AD={5*width_7*LAMBDA} PD={10*LAMBDA+2*width_7}
M8      ref     ref     gnd     gnd  CMOSN   W={width_58}   L={length}
+ AS={5*width_58*LAMBDA} PS={10*LAMBDA+2*width_58} AD={5*width_58*LAMBDA} PD={10*LAMBDA+2*width_58}

* .tran 10u 100m
.ac dec 10 1 100Meg

.control
run

plot v(out) 
plot v(inp) 
plot v(inn)
plot v(inp)-v(inn)

print @M6[gm] 

fourier 10k v(inp)-v(inn)
fourier 10k v(out)

plot (db(v(out))-db(v(inp)-v(inn))) 180/PI*phase(v(out)/(v(inp)-v(inn)))

.endc
