* Telescopic
.include TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param length=0.36u

.param width_1234={0.36*71u}
.param width_5678={0.36*160u}
.param width_910={0.36*142u}
.param width_11={0.36*157u}
.param width_12={0.36*79u}

.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
Iref gnd ref 400u
Vb1 b1 gnd 1.4
Vb2 b2 gnd 0.75

* Transient and AC
* vinp inp gnd dc 0.9 ac 0.01m sin(0.9 0.01m 10k 0 0 0) 
* vinn inn gnd dc 0.9 ac -0.01m sin(0.9 -0.01m 10k 0 0 0)

* Slew Rate
vinp inp gnd pulse(1.8 0 -1n 100p 100p 500n 1u)

* Offset
* vinp inp gnd 0.9

Cc d4 k 2p
Rs k inn 1k

M1      d1     inn      d9     gnd  CMOSN   W={width_1234}   L={length}
+ AS={5*width_1234*LAMBDA} PS={10*LAMBDA+2*width_1234} AD={5*width_1234*LAMBDA} PD={10*LAMBDA+2*width_1234}
M2      d2     inp      d9     gnd  CMOSN   W={width_1234}   L={length}
+ AS={5*width_1234*LAMBDA} PS={10*LAMBDA+2*width_1234} AD={5*width_1234*LAMBDA} PD={10*LAMBDA+2*width_1234}
M3      d3     b1       d1    gnd  CMOSN   W={width_1234}   L={length}
+ AS={5*width_1234*LAMBDA} PS={10*LAMBDA+2*width_1234} AD={5*width_1234*LAMBDA} PD={10*LAMBDA+2*width_1234}
M4      d4     b1       d2    gnd  CMOSN   W={width_1234}   L={length}
+ AS={5*width_1234*LAMBDA} PS={10*LAMBDA+2*width_1234} AD={5*width_1234*LAMBDA} PD={10*LAMBDA+2*width_1234}
M5      d3     b2      d5     vdd  CMOSP   W={width_5678}   L={length}
+ AS={5*width_5678*LAMBDA} PS={10*LAMBDA+2*width_5678} AD={5*width_5678*LAMBDA} PD={10*LAMBDA+2*width_5678}
M6      d4     b2      d6     vdd  CMOSP   W={width_5678}   L={length}
+ AS={5*width_5678*LAMBDA} PS={10*LAMBDA+2*width_5678} AD={5*width_5678*LAMBDA} PD={10*LAMBDA+2*width_5678}
M7      d5     d3       vdd    vdd  CMOSP   W={width_5678}   L={length}
+ AS={5*width_5678*LAMBDA} PS={10*LAMBDA+2*width_5678} AD={5*width_5678*LAMBDA} PD={10*LAMBDA+2*width_5678}
M8      d6     d3       vdd    vdd  CMOSP   W={width_5678}   L={length}
+ AS={5*width_5678*LAMBDA} PS={10*LAMBDA+2*width_5678} AD={5*width_5678*LAMBDA} PD={10*LAMBDA+2*width_5678}


M9      d9    ref      gnd    gnd  CMOSN   W={width_910}   L={length}
+ AS={5*width_910*LAMBDA} PS={10*LAMBDA+2*width_910} AD={5*width_910*LAMBDA} PD={10*LAMBDA+2*width_910}
M10      ref     ref     gnd     gnd  CMOSN   W={width_910}   L={length}
+ AS={5*width_910*LAMBDA} PS={10*LAMBDA+2*width_910} AD={5*width_910*LAMBDA} PD={10*LAMBDA+2*width_910}

M11      inn    d4       vdd    vdd  CMOSP   W={width_11}   L={length}
+ AS={5*width_11*LAMBDA} PS={10*LAMBDA+2*width_11} AD={5*width_11*LAMBDA} PD={10*LAMBDA+2*width_11}
M12      inn    ref      gnd     gnd  CMOSN   W={width_12}   L={length}
+ AS={5*width_12*LAMBDA} PS={10*LAMBDA+2*width_12} AD={5*width_12*LAMBDA} PD={10*LAMBDA+2*width_12}

*.tran 1u 1m
*.op
*.ac dec 10 1 500Meg


* Slew rate & Offset
.tran 0.1n 1u

.control
run


plot v(inp) v(inn) deriv(v(inn))
plot v(inp)-v(inn)

fourier 10k v(inp)-v(inn)
fourier 10k v(inn)

plot (db(v(inn))-db(v(inp)))
plot 180/PI*phase(v(inn)/(v(inp)))

plot (db(v(inn))-db(v(inp))) 180/PI*phase(v(inn)/(v(inp)))

* Slew rate
plot v(inp) V(inn)

.endc
