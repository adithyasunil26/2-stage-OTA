* Telescopic
.include TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param length=0.36u

.param width_1234={0.36*71u}
.param width_5678={0.36*142u}
.param width_910={0.36*142u}
.param width_11={0.36*139u}
.param width_12={0.36*79u}

.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
Iref gnd ref 400u
Vb1 b1 gnd 1.4
Vb2 b2 gnd 0.7

*op
*vinp inp gnd 0.9


* Transient and AC
vinp inp gnd dc 0.9 ac 0.85 sin(0.9 0.85 10k 0 0 0) 
* vinn inn gnd dc 0.9 ac -0.01m sin(0.9 -0.01m 10k 0 0 0)

* Slew Rate
*vinp inp gnd pulse(1 0 -1n 100p 100p 500n 1u)

* Offset
*vinp inp gnd 0

Cc k inn 2p
Rs d4 k 1k

.option scale=0.09u

M1000 d4 b1 d2 gnd CMOSN w=284 l=4
+  ad=1420 pd=578 as=2840 ps=1156
M1001 d4 b2 d6 vdd CMOSP w=640 l=4
+  ad=3200 pd=1290 as=6400 ps=2580
M1002 d6 d3 vdd vdd CMOSP w=640 l=4
+  ad=0 pd=0 as=9540 ps=3846
M1003 d3 b1 d1 gnd CMOSN w=284 l=4
+  ad=1420 pd=578 as=2840 ps=1156
M1004 d9 inp d2 gnd CMOSN w=284 l=4
+  ad=5680 pd=2302 as=0 ps=0
M1005 ref ref gnd gnd CMOSN w=568 l=4
+  ad=2840 pd=1146 as=7080 ps=2862
M1006 d3 b2 d5 vdd CMOSP w=640 l=4
+  ad=3200 pd=1290 as=6400 ps=2580
M1007 d9 inn d1 gnd CMOSN w=284 l=4
+  ad=0 pd=0 as=0 ps=0
M1008 d5 d3 vdd vdd CMOSP w=640 l=4
+  ad=0 pd=0 as=0 ps=0
M1009 inn d4 vdd vdd CMOSP w=628 l=4
+  ad=3140 pd=1266 as=0 ps=0
M1010 gnd ref inn gnd CMOSN w=280 l=4
+  ad=0 pd=0 as=1400 ps=570
M1011 d9 ref gnd gnd CMOSN w=568 l=4
+  ad=0 pd=0 as=0 ps=0
C0 d1 d3 0.02fF
C1 inn d4 0.02fF
C2 d6 d5 0.13fF
C3 d9 inn 0.02fF
C4 b1 d3 0.10fF
C5 inn d3 0.02fF
C6 d6 b2 0.10fF
C7 d6 d3 0.15fF
C8 ref inn 0.03fF
C9 d5 d3 0.12fF
C10 d2 inn 0.09fF
C11 vdd inn 0.02fF
C12 d9 inp 0.10fF
C13 d4 d3 0.14fF
C14 d1 inn 0.11fF
C15 vdd d6 0.04fF
C16 b2 d3 0.21fF
C17 gnd d4 0.02fF
C18 vdd d5 0.06fF
C19 d9 ref 0.23fF
C20 gnd d9 0.04fF
C21 d2 d4 0.02fF
C22 vdd d4 0.21fF
C23 gnd b2 0.16fF
C24 d9 d2 0.02fF
C25 gnd inp 0.08fF
C26 d1 d4 0.02fF
C27 vdd b2 0.23fF
C28 gnd d3 0.16fF
C29 gnd inn 0.08fF
C30 b1 d4 0.21fF
C31 vdd d3 0.35fF
C32 gnd ref 0.04fF
C33 d9 gnd 0.06fF
C34 inp gnd 0.13fF
C35 inn gnd 0.13fF
C36 ref gnd 0.49fF
C37 d2 gnd 0.06fF
C38 d1 gnd 0.06fF
C39 b1 gnd 0.04fF
C40 inn gnd 0.91fF
C41 d6 gnd 0.00fF
C42 d5 gnd 0.00fF
C43 d4 gnd 0.07fF
C44 b2 gnd 0.04fF
C45 d3 gnd 0.09fF
C46 gnd gnd 15.36fF
C47 vdd gnd 70.82fF


.tran 1u 1m
*.op
*.ac dec 10 1 1000Meg
*.dc vinp 0 1.8 0.01


* Slew rate & Offset
*.tran 0.01u 1u

.control
run
set hcopypscolor = 1
set color0=white
set color1=black

*plot v(inp) v(inn) deriv(v(inn))
*plot v(inp)-v(inn)

*fourier 10k v(inp)-v(inn)
fourier 10k v(inn)

*plot (db(v(inn))-db(v(inp)))
*plot 180/PI*phase(v(inn)/(v(inp)))

*plot (db(v(inn))-db(v(inp))) 180/PI*phase(v(inn)/(v(inp)))


* Slew rate
plot v(inp) V(inn)
*plot deriv(v(inn))

*plot v(inn)
*plot deriv(v(inn))
.endc
