magic
tech scmos
timestamp 1638481995
<< nwell >>
rect -6 -6 100 586
<< ntransistor >>
rect 119 280 123 564
rect 139 280 143 564
rect 119 -19 123 265
rect 139 -19 143 265
rect 159 -19 163 297
rect 179 -19 183 549
rect 199 -19 203 549
<< ptransistor >>
rect 5 0 9 568
rect 25 0 29 568
rect 45 0 49 568
rect 65 0 69 568
rect 85 12 89 568
<< ndiffusion >>
rect 114 284 119 564
rect 118 280 119 284
rect 123 535 128 564
rect 123 531 124 535
rect 123 280 128 531
rect 134 284 139 564
rect 138 280 139 284
rect 143 520 148 564
rect 143 516 144 520
rect 143 280 148 516
rect 158 293 159 297
rect 118 261 119 265
rect 114 -19 119 261
rect 123 68 128 265
rect 123 64 124 68
rect 123 -19 128 64
rect 138 261 139 265
rect 134 -19 139 261
rect 143 68 148 265
rect 143 64 144 68
rect 143 -19 148 64
rect 154 -19 159 293
rect 163 -15 168 297
rect 163 -19 164 -15
rect 174 -15 179 549
rect 178 -19 179 -15
rect 183 68 188 549
rect 183 64 184 68
rect 183 -19 188 64
rect 194 -15 199 549
rect 198 -19 199 -15
rect 203 545 204 549
rect 203 304 208 545
rect 203 300 204 304
rect 203 -19 208 300
<< pdiffusion >>
rect 4 564 5 568
rect 0 0 5 564
rect 9 556 14 568
rect 9 552 10 556
rect 9 0 14 552
rect 24 564 25 568
rect 20 0 25 564
rect 29 546 34 568
rect 29 542 30 546
rect 29 0 34 542
rect 40 556 45 568
rect 44 552 45 556
rect 40 0 45 552
rect 49 535 54 568
rect 49 531 50 535
rect 49 14 54 531
rect 49 10 50 14
rect 49 0 54 10
rect 60 546 65 568
rect 64 542 65 546
rect 60 0 65 542
rect 69 520 74 568
rect 69 516 70 520
rect 69 9 74 516
rect 84 564 85 568
rect 80 12 85 564
rect 89 274 94 568
rect 89 270 90 274
rect 89 12 94 270
rect 69 5 70 9
rect 69 0 74 5
<< ndcontact >>
rect 114 280 118 284
rect 124 531 128 535
rect 134 280 138 284
rect 144 516 148 520
rect 154 293 158 297
rect 114 261 118 265
rect 124 64 128 68
rect 134 261 138 265
rect 144 64 148 68
rect 164 -19 168 -15
rect 174 -19 178 -15
rect 184 64 188 68
rect 194 -19 198 -15
rect 204 545 208 549
rect 204 300 208 304
<< pdcontact >>
rect 0 564 4 568
rect 10 552 14 556
rect 20 564 24 568
rect 30 542 34 546
rect 40 552 44 556
rect 50 531 54 535
rect 50 10 54 14
rect 60 542 64 546
rect 70 516 74 520
rect 80 564 84 568
rect 90 270 94 274
rect 70 5 74 9
<< psubstratepcontact >>
rect 114 -38 118 -34
rect 124 -38 128 -34
rect 134 -38 138 -34
rect 144 -38 148 -34
rect 154 -38 158 -34
rect 164 -38 168 -34
rect 174 -38 178 -34
rect 184 -38 188 -34
rect 194 -38 198 -34
rect 204 -38 208 -34
<< nsubstratencontact >>
rect 0 578 4 582
rect 10 578 14 582
rect 20 578 24 582
rect 30 578 34 582
rect 40 578 44 582
rect 50 578 54 582
rect 60 578 64 582
rect 70 578 74 582
rect 80 578 84 582
rect 90 578 94 582
<< polysilicon >>
rect 5 568 9 571
rect 25 568 29 571
rect 45 568 49 571
rect 65 568 69 571
rect 85 568 89 571
rect 119 564 123 567
rect 139 564 143 567
rect 179 549 183 552
rect 199 549 203 552
rect 159 297 163 300
rect 119 277 123 280
rect 139 277 143 280
rect 119 265 123 268
rect 139 265 143 268
rect 85 9 89 12
rect 5 -2 9 0
rect 25 -2 29 0
rect 45 -2 49 0
rect 65 -2 69 0
rect 119 -22 123 -19
rect 139 -22 143 -19
rect 159 -22 163 -19
rect 179 -22 183 -19
rect 199 -22 203 -19
<< polycontact >>
rect 119 567 123 571
rect 139 567 143 571
rect 179 552 183 556
rect 199 552 203 556
rect 159 300 163 304
rect 85 5 89 9
rect 5 -6 9 -2
rect 25 -6 29 -2
rect 45 -6 49 -2
rect 65 -6 69 -2
rect 119 -26 123 -22
rect 139 -26 143 -22
<< metal1 >>
rect -6 582 100 586
rect -6 578 0 582
rect 4 578 10 582
rect 14 578 20 582
rect 24 578 30 582
rect 34 578 40 582
rect 44 578 50 582
rect 54 578 60 582
rect 64 578 70 582
rect 74 578 80 582
rect 84 578 90 582
rect 94 578 100 582
rect -6 574 100 578
rect 0 568 4 574
rect 20 568 24 574
rect 80 568 84 574
rect 123 567 139 571
rect 14 552 40 556
rect 183 552 199 556
rect 203 552 208 556
rect 204 549 208 552
rect 34 542 60 546
rect 54 531 124 535
rect 74 516 144 520
rect 150 308 154 312
rect 150 293 154 303
rect 163 300 204 304
rect 94 270 102 274
rect 114 265 118 280
rect 134 265 138 280
rect 128 64 144 68
rect 148 64 184 68
rect 25 10 50 14
rect 25 -2 29 10
rect 74 5 85 9
rect 9 -6 25 -2
rect 49 -6 65 -2
rect 115 -26 119 -22
rect 135 -26 139 -22
rect 164 -30 168 -19
rect 174 -30 178 -19
rect 194 -30 198 -19
rect 108 -34 214 -30
rect 108 -38 114 -34
rect 118 -38 124 -34
rect 128 -38 134 -34
rect 138 -38 144 -34
rect 148 -38 154 -34
rect 158 -38 164 -34
rect 168 -38 174 -34
rect 178 -38 184 -34
rect 188 -38 194 -34
rect 198 -38 204 -34
rect 208 -38 214 -34
rect 108 -42 214 -38
<< m2contact >>
rect 149 303 154 308
rect 102 269 107 274
<< metal2 >>
rect 149 274 153 303
rect 107 270 153 274
<< labels >>
rlabel metal1 56 -5 56 -5 1 b2
rlabel metal1 82 571 82 571 1 vdd!
rlabel metal1 104 518 104 518 1 d4
rlabel metal1 104 533 104 533 1 d3
rlabel metal1 36 554 36 554 1 d5
rlabel metal1 57 544 57 544 1 d6
rlabel metal1 131 568 131 568 1 b1
rlabel metal1 190 554 190 554 1 ref
rlabel metal1 152 310 152 310 1 out
rlabel metal1 137 -24 137 -24 1 inp
rlabel metal1 117 -24 117 -24 1 inn
rlabel metal1 151 66 151 66 1 d9
rlabel metal1 116 266 116 266 1 d1
rlabel metal1 136 267 136 267 1 d2
rlabel metal1 196 -25 196 -25 1 gnd!
<< end >>
