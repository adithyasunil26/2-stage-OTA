magic
tech scmos
timestamp 1638491757
<< nwell >>
rect -6 -6 100 586
<< ntransistor >>
rect 119 280 123 564
rect 139 280 143 564
rect 119 -19 123 265
rect 139 -19 143 265
rect 159 -19 163 297
rect 179 -19 183 549
rect 199 -19 203 549
<< ptransistor >>
rect 5 0 9 568
rect 25 0 29 568
rect 45 0 49 568
rect 65 0 69 568
rect 85 12 89 568
<< ndiffusion >>
rect 114 284 119 564
rect 118 280 119 284
rect 123 535 128 564
rect 123 531 124 535
rect 123 280 128 531
rect 134 284 139 564
rect 138 280 139 284
rect 143 520 148 564
rect 143 516 144 520
rect 143 280 148 516
rect 158 293 159 297
rect 118 261 119 265
rect 114 -19 119 261
rect 123 68 128 265
rect 123 64 124 68
rect 123 -19 128 64
rect 138 261 139 265
rect 134 -19 139 261
rect 143 68 148 265
rect 143 64 144 68
rect 143 -19 148 64
rect 154 -19 159 293
rect 163 -15 168 297
rect 163 -19 164 -15
rect 174 -15 179 549
rect 178 -19 179 -15
rect 183 68 188 549
rect 183 64 184 68
rect 183 -19 188 64
rect 194 -15 199 549
rect 198 -19 199 -15
rect 203 545 204 549
rect 203 304 208 545
rect 203 300 204 304
rect 203 -19 208 300
<< pdiffusion >>
rect 4 564 5 568
rect 0 0 5 564
rect 9 556 14 568
rect 9 552 10 556
rect 9 0 14 552
rect 24 564 25 568
rect 20 0 25 564
rect 29 546 34 568
rect 29 542 30 546
rect 29 0 34 542
rect 40 556 45 568
rect 44 552 45 556
rect 40 0 45 552
rect 49 535 54 568
rect 49 531 50 535
rect 49 14 54 531
rect 49 10 50 14
rect 49 0 54 10
rect 60 546 65 568
rect 64 542 65 546
rect 60 0 65 542
rect 69 520 74 568
rect 69 516 70 520
rect 69 9 74 516
rect 84 564 85 568
rect 80 12 85 564
rect 89 274 94 568
rect 89 270 90 274
rect 89 12 94 270
rect 69 5 70 9
rect 69 0 74 5
<< ndcontact >>
rect 114 280 118 284
rect 124 531 128 535
rect 134 280 138 284
rect 144 516 148 520
rect 154 293 158 297
rect 114 261 118 265
rect 124 64 128 68
rect 134 261 138 265
rect 144 64 148 68
rect 164 -19 168 -15
rect 174 -19 178 -15
rect 184 64 188 68
rect 194 -19 198 -15
rect 204 545 208 549
rect 204 300 208 304
<< pdcontact >>
rect 0 564 4 568
rect 10 552 14 556
rect 20 564 24 568
rect 30 542 34 546
rect 40 552 44 556
rect 50 531 54 535
rect 50 10 54 14
rect 60 542 64 546
rect 70 516 74 520
rect 80 564 84 568
rect 90 270 94 274
rect 70 5 74 9
<< psubstratepcontact >>
rect -26 602 -22 606
rect -16 602 -12 606
rect -6 602 -2 606
rect 4 602 8 606
rect 14 602 18 606
rect 24 602 28 606
rect 34 602 38 606
rect 44 602 48 606
rect 54 602 58 606
rect 64 602 68 606
rect 74 602 78 606
rect 84 602 88 606
rect 94 602 98 606
rect 104 602 108 606
rect 114 602 118 606
rect 124 602 128 606
rect 134 602 138 606
rect 144 602 148 606
rect 154 602 158 606
rect 164 602 168 606
rect 174 602 178 606
rect 184 602 188 606
rect 194 602 198 606
rect 204 602 208 606
rect 214 602 218 606
rect 224 602 228 606
rect -26 592 -22 596
rect 224 592 228 596
rect -26 582 -22 586
rect 114 583 118 587
rect 124 583 128 587
rect 134 583 138 587
rect 144 583 148 587
rect 154 583 158 587
rect 164 583 168 587
rect 174 583 178 587
rect 184 583 188 587
rect 194 583 198 587
rect 204 583 208 587
rect 214 583 218 587
rect 224 582 228 586
rect -26 572 -22 576
rect 159 572 163 576
rect 224 572 228 576
rect -26 562 -22 566
rect -26 552 -22 556
rect -26 542 -22 546
rect -26 532 -22 536
rect -26 522 -22 526
rect -26 512 -22 516
rect -26 502 -22 506
rect -26 492 -22 496
rect -26 482 -22 486
rect -26 472 -22 476
rect -26 462 -22 466
rect -26 452 -22 456
rect -26 442 -22 446
rect -26 432 -22 436
rect -26 422 -22 426
rect -26 412 -22 416
rect -26 402 -22 406
rect -26 392 -22 396
rect -26 382 -22 386
rect -26 372 -22 376
rect -26 362 -22 366
rect -26 352 -22 356
rect -26 342 -22 346
rect -26 332 -22 336
rect -26 322 -22 326
rect -26 312 -22 316
rect -26 302 -22 306
rect -26 292 -22 296
rect -26 282 -22 286
rect -26 272 -22 276
rect -26 262 -22 266
rect -26 252 -22 256
rect -26 242 -22 246
rect -26 232 -22 236
rect -26 222 -22 226
rect -26 212 -22 216
rect -26 202 -22 206
rect -26 192 -22 196
rect -26 182 -22 186
rect -26 172 -22 176
rect -26 162 -22 166
rect -26 152 -22 156
rect -26 142 -22 146
rect -26 132 -22 136
rect -26 122 -22 126
rect -26 112 -22 116
rect -26 102 -22 106
rect -26 92 -22 96
rect -26 82 -22 86
rect -26 72 -22 76
rect -26 62 -22 66
rect -26 52 -22 56
rect -26 42 -22 46
rect -26 32 -22 36
rect -26 22 -22 26
rect -26 12 -22 16
rect -26 2 -22 6
rect 159 562 163 566
rect 224 562 228 566
rect 159 552 163 556
rect 224 552 228 556
rect 159 542 163 546
rect 159 532 163 536
rect 159 522 163 526
rect 159 512 163 516
rect 159 502 163 506
rect 159 492 163 496
rect 159 482 163 486
rect 159 472 163 476
rect 159 462 163 466
rect 159 452 163 456
rect 159 442 163 446
rect 159 432 163 436
rect 159 422 163 426
rect 159 412 163 416
rect 159 402 163 406
rect 159 392 163 396
rect 159 382 163 386
rect 159 372 163 376
rect 159 362 163 366
rect 159 352 163 356
rect 159 342 163 346
rect 159 332 163 336
rect -26 -8 -22 -4
rect -26 -18 -22 -14
rect -16 -19 -12 -15
rect -6 -19 -2 -15
rect 4 -19 8 -15
rect 14 -19 18 -15
rect 24 -19 28 -15
rect 34 -19 38 -15
rect 44 -19 48 -15
rect 54 -19 58 -15
rect 64 -19 68 -15
rect 74 -19 78 -15
rect 84 -19 88 -15
rect 94 -19 98 -15
rect 224 542 228 546
rect 224 532 228 536
rect 224 522 228 526
rect 224 512 228 516
rect 224 502 228 506
rect 224 492 228 496
rect 224 482 228 486
rect 224 472 228 476
rect 224 462 228 466
rect 224 452 228 456
rect 224 442 228 446
rect 224 432 228 436
rect 224 422 228 426
rect 224 412 228 416
rect 224 402 228 406
rect 224 392 228 396
rect 224 382 228 386
rect 224 372 228 376
rect 224 362 228 366
rect 224 352 228 356
rect 224 342 228 346
rect 224 332 228 336
rect 224 322 228 326
rect 224 312 228 316
rect 224 302 228 306
rect 224 292 228 296
rect 224 282 228 286
rect 224 272 228 276
rect 224 262 228 266
rect 224 252 228 256
rect 224 242 228 246
rect 224 232 228 236
rect 224 222 228 226
rect 224 212 228 216
rect 224 202 228 206
rect 224 192 228 196
rect 224 182 228 186
rect 224 172 228 176
rect 224 162 228 166
rect 224 152 228 156
rect 224 142 228 146
rect 224 132 228 136
rect 224 122 228 126
rect 224 112 228 116
rect 224 102 228 106
rect 224 92 228 96
rect 224 82 228 86
rect 224 72 228 76
rect 224 62 228 66
rect 224 52 228 56
rect 224 42 228 46
rect 224 32 228 36
rect 224 22 228 26
rect 224 12 228 16
rect 224 2 228 6
rect 224 -8 228 -4
rect 224 -18 228 -14
rect -26 -28 -22 -24
rect 224 -28 228 -24
rect -26 -38 -22 -34
rect -16 -38 -12 -34
rect -6 -38 -2 -34
rect 4 -38 8 -34
rect 14 -38 18 -34
rect 24 -38 28 -34
rect 34 -38 38 -34
rect 44 -38 48 -34
rect 54 -38 58 -34
rect 64 -38 68 -34
rect 74 -38 78 -34
rect 84 -38 88 -34
rect 94 -38 98 -34
rect 104 -38 108 -34
rect 114 -38 118 -34
rect 124 -38 128 -34
rect 134 -38 138 -34
rect 144 -38 148 -34
rect 154 -38 158 -34
rect 164 -38 168 -34
rect 174 -38 178 -34
rect 184 -38 188 -34
rect 194 -38 198 -34
rect 204 -38 208 -34
rect 214 -38 218 -34
rect 224 -38 228 -34
<< nsubstratencontact >>
rect 0 578 4 582
rect 10 578 14 582
rect 20 578 24 582
rect 30 578 34 582
rect 40 578 44 582
rect 50 578 54 582
rect 60 578 64 582
rect 70 578 74 582
rect 80 578 84 582
rect 90 578 94 582
<< polysilicon >>
rect 5 568 9 571
rect 25 568 29 571
rect 45 568 49 571
rect 65 568 69 571
rect 85 568 89 571
rect 119 564 123 567
rect 139 564 143 567
rect 179 549 183 552
rect 199 549 203 552
rect 159 297 163 300
rect 119 277 123 280
rect 139 277 143 280
rect 119 265 123 268
rect 139 265 143 268
rect 85 9 89 12
rect 5 -2 9 0
rect 25 -2 29 0
rect 45 -2 49 0
rect 65 -2 69 0
rect 119 -22 123 -19
rect 139 -22 143 -19
rect 159 -22 163 -19
rect 179 -22 183 -19
rect 199 -22 203 -19
<< polycontact >>
rect 119 567 123 571
rect 139 567 143 571
rect 179 552 183 556
rect 199 552 203 556
rect 159 300 163 304
rect 85 5 89 9
rect 5 -6 9 -2
rect 25 -6 29 -2
rect 45 -6 49 -2
rect 65 -6 69 -2
rect 119 -26 123 -22
rect 139 -26 143 -22
<< metal1 >>
rect -30 606 232 610
rect -30 602 -26 606
rect -22 602 -16 606
rect -12 602 -6 606
rect -2 602 4 606
rect 8 602 14 606
rect 18 602 24 606
rect 28 602 34 606
rect 38 602 44 606
rect 48 602 54 606
rect 58 602 64 606
rect 68 602 74 606
rect 78 602 84 606
rect 88 602 94 606
rect 98 602 104 606
rect 108 602 114 606
rect 118 602 124 606
rect 128 602 134 606
rect 138 602 144 606
rect 148 602 154 606
rect 158 602 164 606
rect 168 602 174 606
rect 178 602 184 606
rect 188 602 194 606
rect 198 602 204 606
rect 208 602 214 606
rect 218 602 224 606
rect 228 602 232 606
rect -30 598 232 602
rect -30 596 -18 598
rect -30 592 -26 596
rect -22 592 -18 596
rect -30 586 -18 592
rect 220 596 232 598
rect 220 592 224 596
rect 228 592 232 596
rect 220 591 232 592
rect 108 587 232 591
rect -30 582 -26 586
rect -22 582 -18 586
rect -30 576 -18 582
rect -30 572 -26 576
rect -22 572 -18 576
rect -6 582 100 586
rect -6 578 0 582
rect 4 578 10 582
rect 14 578 20 582
rect 24 578 30 582
rect 34 578 40 582
rect 44 578 50 582
rect 54 578 60 582
rect 64 578 70 582
rect 74 578 80 582
rect 84 578 90 582
rect 94 578 100 582
rect 108 583 114 587
rect 118 583 124 587
rect 128 583 134 587
rect 138 583 144 587
rect 148 583 154 587
rect 158 583 164 587
rect 168 583 174 587
rect 178 583 184 587
rect 188 583 194 587
rect 198 583 204 587
rect 208 583 214 587
rect 218 586 232 587
rect 218 583 224 586
rect 108 582 224 583
rect 228 582 232 586
rect 108 579 232 582
rect -6 574 100 578
rect 155 576 167 579
rect -30 566 -18 572
rect -30 562 -26 566
rect -22 562 -18 566
rect 0 568 4 574
rect 20 568 24 574
rect 80 568 84 574
rect 155 572 159 576
rect 163 572 167 576
rect 123 567 139 571
rect 155 566 167 572
rect -30 556 -18 562
rect 155 562 159 566
rect 163 562 167 566
rect 155 556 167 562
rect 220 576 232 579
rect 220 572 224 576
rect 228 572 232 576
rect 220 566 232 572
rect 220 562 224 566
rect 228 562 232 566
rect 220 556 232 562
rect -30 552 -26 556
rect -22 552 -18 556
rect 14 552 40 556
rect 155 552 159 556
rect 163 552 167 556
rect 183 552 199 556
rect 203 552 208 556
rect -30 546 -18 552
rect 155 546 167 552
rect -30 542 -26 546
rect -22 542 -18 546
rect 34 542 60 546
rect 155 542 159 546
rect 163 542 167 546
rect 204 549 208 552
rect 220 552 224 556
rect 228 552 232 556
rect 220 546 232 552
rect -30 536 -18 542
rect -30 532 -26 536
rect -22 532 -18 536
rect 155 536 167 542
rect -30 526 -18 532
rect 54 531 124 535
rect 155 532 159 536
rect 163 532 167 536
rect -30 522 -26 526
rect -22 522 -18 526
rect -30 516 -18 522
rect 155 526 167 532
rect 155 522 159 526
rect 163 522 167 526
rect 74 516 144 520
rect 155 516 167 522
rect -30 512 -26 516
rect -22 512 -18 516
rect -30 506 -18 512
rect -30 502 -26 506
rect -22 502 -18 506
rect -30 496 -18 502
rect -30 492 -26 496
rect -22 492 -18 496
rect -30 486 -18 492
rect -30 482 -26 486
rect -22 482 -18 486
rect -30 476 -18 482
rect -30 472 -26 476
rect -22 472 -18 476
rect -30 466 -18 472
rect -30 462 -26 466
rect -22 462 -18 466
rect -30 456 -18 462
rect -30 452 -26 456
rect -22 452 -18 456
rect -30 446 -18 452
rect -30 442 -26 446
rect -22 442 -18 446
rect -30 436 -18 442
rect -30 432 -26 436
rect -22 432 -18 436
rect -30 426 -18 432
rect -30 422 -26 426
rect -22 422 -18 426
rect -30 416 -18 422
rect -30 412 -26 416
rect -22 412 -18 416
rect -30 406 -18 412
rect -30 402 -26 406
rect -22 402 -18 406
rect -30 396 -18 402
rect -30 392 -26 396
rect -22 392 -18 396
rect -30 386 -18 392
rect -30 382 -26 386
rect -22 382 -18 386
rect -30 376 -18 382
rect -30 372 -26 376
rect -22 372 -18 376
rect -30 366 -18 372
rect -30 362 -26 366
rect -22 362 -18 366
rect -30 356 -18 362
rect -30 352 -26 356
rect -22 352 -18 356
rect -30 346 -18 352
rect -30 342 -26 346
rect -22 342 -18 346
rect -30 336 -18 342
rect -30 332 -26 336
rect -22 332 -18 336
rect -30 326 -18 332
rect 155 512 159 516
rect 163 512 167 516
rect 155 506 167 512
rect 155 502 159 506
rect 163 502 167 506
rect 155 496 167 502
rect 155 492 159 496
rect 163 492 167 496
rect 155 486 167 492
rect 155 482 159 486
rect 163 482 167 486
rect 155 476 167 482
rect 155 472 159 476
rect 163 472 167 476
rect 155 466 167 472
rect 155 462 159 466
rect 163 462 167 466
rect 155 456 167 462
rect 155 452 159 456
rect 163 452 167 456
rect 155 446 167 452
rect 155 442 159 446
rect 163 442 167 446
rect 155 436 167 442
rect 155 432 159 436
rect 163 432 167 436
rect 155 426 167 432
rect 155 422 159 426
rect 163 422 167 426
rect 155 416 167 422
rect 155 412 159 416
rect 163 412 167 416
rect 155 406 167 412
rect 155 402 159 406
rect 163 402 167 406
rect 155 396 167 402
rect 155 392 159 396
rect 163 392 167 396
rect 155 386 167 392
rect 155 382 159 386
rect 163 382 167 386
rect 155 376 167 382
rect 155 372 159 376
rect 163 372 167 376
rect 155 366 167 372
rect 155 362 159 366
rect 163 362 167 366
rect 155 356 167 362
rect 155 352 159 356
rect 163 352 167 356
rect 155 346 167 352
rect 155 342 159 346
rect 163 342 167 346
rect 155 336 167 342
rect 155 332 159 336
rect 163 332 167 336
rect 155 326 167 332
rect 220 542 224 546
rect 228 542 232 546
rect 220 536 232 542
rect 220 532 224 536
rect 228 532 232 536
rect 220 526 232 532
rect 220 522 224 526
rect 228 522 232 526
rect 220 516 232 522
rect 220 512 224 516
rect 228 512 232 516
rect 220 506 232 512
rect 220 502 224 506
rect 228 502 232 506
rect 220 496 232 502
rect 220 492 224 496
rect 228 492 232 496
rect 220 486 232 492
rect 220 482 224 486
rect 228 482 232 486
rect 220 476 232 482
rect 220 472 224 476
rect 228 472 232 476
rect 220 466 232 472
rect 220 462 224 466
rect 228 462 232 466
rect 220 456 232 462
rect 220 452 224 456
rect 228 452 232 456
rect 220 446 232 452
rect 220 442 224 446
rect 228 442 232 446
rect 220 436 232 442
rect 220 432 224 436
rect 228 432 232 436
rect 220 426 232 432
rect 220 422 224 426
rect 228 422 232 426
rect 220 416 232 422
rect 220 412 224 416
rect 228 412 232 416
rect 220 406 232 412
rect 220 402 224 406
rect 228 402 232 406
rect 220 396 232 402
rect 220 392 224 396
rect 228 392 232 396
rect 220 386 232 392
rect 220 382 224 386
rect 228 382 232 386
rect 220 376 232 382
rect 220 372 224 376
rect 228 372 232 376
rect 220 366 232 372
rect 220 362 224 366
rect 228 362 232 366
rect 220 356 232 362
rect 220 352 224 356
rect 228 352 232 356
rect 220 346 232 352
rect 220 342 224 346
rect 228 342 232 346
rect 220 336 232 342
rect 220 332 224 336
rect 228 332 232 336
rect 220 326 232 332
rect -30 322 -26 326
rect -22 322 -18 326
rect -30 316 -18 322
rect -30 312 -26 316
rect -22 312 -18 316
rect 220 322 224 326
rect 228 322 232 326
rect 220 316 232 322
rect 220 312 224 316
rect 228 312 232 316
rect -30 306 -18 312
rect 150 308 154 312
rect -30 302 -26 306
rect -22 302 -18 306
rect 220 306 232 312
rect -30 296 -18 302
rect -30 292 -26 296
rect -22 292 -18 296
rect 150 293 154 303
rect 163 300 204 304
rect 220 302 224 306
rect 228 302 232 306
rect 220 296 232 302
rect -30 286 -18 292
rect -30 282 -26 286
rect -22 282 -18 286
rect 220 292 224 296
rect 228 292 232 296
rect 220 286 232 292
rect -30 276 -18 282
rect -30 272 -26 276
rect -22 272 -18 276
rect -30 266 -18 272
rect 94 270 102 274
rect -30 262 -26 266
rect -22 262 -18 266
rect -30 256 -18 262
rect 114 265 118 280
rect 134 265 138 280
rect 220 282 224 286
rect 228 282 232 286
rect 220 276 232 282
rect 220 272 224 276
rect 228 272 232 276
rect 220 266 232 272
rect 220 262 224 266
rect 228 262 232 266
rect -30 252 -26 256
rect -22 252 -18 256
rect -30 246 -18 252
rect -30 242 -26 246
rect -22 242 -18 246
rect -30 236 -18 242
rect -30 232 -26 236
rect -22 232 -18 236
rect -30 226 -18 232
rect -30 222 -26 226
rect -22 222 -18 226
rect -30 216 -18 222
rect -30 212 -26 216
rect -22 212 -18 216
rect -30 206 -18 212
rect -30 202 -26 206
rect -22 202 -18 206
rect -30 196 -18 202
rect -30 192 -26 196
rect -22 192 -18 196
rect -30 186 -18 192
rect -30 182 -26 186
rect -22 182 -18 186
rect -30 176 -18 182
rect -30 172 -26 176
rect -22 172 -18 176
rect -30 166 -18 172
rect -30 162 -26 166
rect -22 162 -18 166
rect -30 156 -18 162
rect -30 152 -26 156
rect -22 152 -18 156
rect -30 146 -18 152
rect -30 142 -26 146
rect -22 142 -18 146
rect -30 136 -18 142
rect -30 132 -26 136
rect -22 132 -18 136
rect -30 126 -18 132
rect -30 122 -26 126
rect -22 122 -18 126
rect -30 116 -18 122
rect -30 112 -26 116
rect -22 112 -18 116
rect -30 106 -18 112
rect -30 102 -26 106
rect -22 102 -18 106
rect -30 96 -18 102
rect -30 92 -26 96
rect -22 92 -18 96
rect -30 86 -18 92
rect -30 82 -26 86
rect -22 82 -18 86
rect -30 76 -18 82
rect -30 72 -26 76
rect -22 72 -18 76
rect -30 66 -18 72
rect 220 256 232 262
rect 220 252 224 256
rect 228 252 232 256
rect 220 246 232 252
rect 220 242 224 246
rect 228 242 232 246
rect 220 236 232 242
rect 220 232 224 236
rect 228 232 232 236
rect 220 226 232 232
rect 220 222 224 226
rect 228 222 232 226
rect 220 216 232 222
rect 220 212 224 216
rect 228 212 232 216
rect 220 206 232 212
rect 220 202 224 206
rect 228 202 232 206
rect 220 196 232 202
rect 220 192 224 196
rect 228 192 232 196
rect 220 186 232 192
rect 220 182 224 186
rect 228 182 232 186
rect 220 176 232 182
rect 220 172 224 176
rect 228 172 232 176
rect 220 166 232 172
rect 220 162 224 166
rect 228 162 232 166
rect 220 156 232 162
rect 220 152 224 156
rect 228 152 232 156
rect 220 146 232 152
rect 220 142 224 146
rect 228 142 232 146
rect 220 136 232 142
rect 220 132 224 136
rect 228 132 232 136
rect 220 126 232 132
rect 220 122 224 126
rect 228 122 232 126
rect 220 116 232 122
rect 220 112 224 116
rect 228 112 232 116
rect 220 106 232 112
rect 220 102 224 106
rect 228 102 232 106
rect 220 96 232 102
rect 220 92 224 96
rect 228 92 232 96
rect 220 86 232 92
rect 220 82 224 86
rect 228 82 232 86
rect 220 76 232 82
rect 220 72 224 76
rect 228 72 232 76
rect -30 62 -26 66
rect -22 62 -18 66
rect 128 64 144 68
rect 148 64 184 68
rect 220 66 232 72
rect -30 56 -18 62
rect -30 52 -26 56
rect -22 52 -18 56
rect -30 46 -18 52
rect -30 42 -26 46
rect -22 42 -18 46
rect -30 36 -18 42
rect -30 32 -26 36
rect -22 32 -18 36
rect -30 26 -18 32
rect -30 22 -26 26
rect -22 22 -18 26
rect -30 16 -18 22
rect -30 12 -26 16
rect -22 12 -18 16
rect 220 62 224 66
rect 228 62 232 66
rect 220 56 232 62
rect 220 52 224 56
rect 228 52 232 56
rect 220 46 232 52
rect 220 42 224 46
rect 228 42 232 46
rect 220 36 232 42
rect 220 32 224 36
rect 228 32 232 36
rect 220 26 232 32
rect 220 22 224 26
rect 228 22 232 26
rect 220 16 232 22
rect -30 6 -18 12
rect -30 2 -26 6
rect -22 2 -18 6
rect -30 -4 -18 2
rect 25 10 50 14
rect 220 12 224 16
rect 228 12 232 16
rect 25 -2 29 10
rect 74 5 85 9
rect 220 6 232 12
rect 220 2 224 6
rect 228 2 232 6
rect -30 -8 -26 -4
rect -22 -8 -18 -4
rect 9 -6 25 -2
rect 49 -6 65 -2
rect 220 -4 232 2
rect -30 -12 -18 -8
rect 220 -8 224 -4
rect 228 -8 232 -4
rect -30 -14 103 -12
rect -30 -18 -26 -14
rect -22 -15 103 -14
rect 220 -14 232 -8
rect -22 -18 -16 -15
rect -30 -19 -16 -18
rect -12 -19 -6 -15
rect -2 -19 4 -15
rect 8 -19 14 -15
rect 18 -19 24 -15
rect 28 -19 34 -15
rect 38 -19 44 -15
rect 48 -19 54 -15
rect 58 -19 64 -15
rect 68 -19 74 -15
rect 78 -19 84 -15
rect 88 -19 94 -15
rect 98 -19 103 -15
rect -30 -22 103 -19
rect -30 -24 -18 -22
rect -30 -28 -26 -24
rect -22 -28 -18 -24
rect 115 -26 119 -22
rect 135 -26 139 -22
rect -30 -30 -18 -28
rect 164 -30 168 -19
rect 174 -30 178 -19
rect 194 -30 198 -19
rect 220 -18 224 -14
rect 228 -18 232 -14
rect 220 -24 232 -18
rect 220 -28 224 -24
rect 228 -28 232 -24
rect 220 -30 232 -28
rect -30 -34 232 -30
rect -30 -38 -26 -34
rect -22 -38 -16 -34
rect -12 -38 -6 -34
rect -2 -38 4 -34
rect 8 -38 14 -34
rect 18 -38 24 -34
rect 28 -38 34 -34
rect 38 -38 44 -34
rect 48 -38 54 -34
rect 58 -38 64 -34
rect 68 -38 74 -34
rect 78 -38 84 -34
rect 88 -38 94 -34
rect 98 -38 104 -34
rect 108 -38 114 -34
rect 118 -38 124 -34
rect 128 -38 134 -34
rect 138 -38 144 -34
rect 148 -38 154 -34
rect 158 -38 164 -34
rect 168 -38 174 -34
rect 178 -38 184 -34
rect 188 -38 194 -34
rect 198 -38 204 -34
rect 208 -38 214 -34
rect 218 -38 224 -34
rect 228 -38 232 -34
rect -30 -42 232 -38
<< m2contact >>
rect 149 303 154 308
rect 102 269 107 274
<< metal2 >>
rect 149 274 153 303
rect 107 270 153 274
<< labels >>
rlabel metal1 56 -5 56 -5 1 b2
rlabel metal1 82 571 82 571 1 vdd!
rlabel metal1 104 518 104 518 1 d4
rlabel metal1 104 533 104 533 1 d3
rlabel metal1 36 554 36 554 1 d5
rlabel metal1 57 544 57 544 1 d6
rlabel metal1 131 568 131 568 1 b1
rlabel metal1 190 554 190 554 1 ref
rlabel metal1 152 310 152 310 1 out
rlabel metal1 137 -24 137 -24 1 inp
rlabel metal1 117 -24 117 -24 1 inn
rlabel metal1 151 66 151 66 1 d9
rlabel metal1 116 266 116 266 1 d1
rlabel metal1 136 267 136 267 1 d2
rlabel metal1 196 -25 196 -25 1 gnd!
<< end >>
