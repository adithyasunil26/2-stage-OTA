magic
tech scmos
timestamp 1638698369
<< nwell >>
rect 6 90 670 196
<< ntransistor >>
rect -7 67 277 71
rect 292 67 576 71
rect -7 47 277 51
rect 292 47 576 51
rect 29 27 309 31
rect -7 7 561 11
rect -7 -13 561 -9
<< ptransistor >>
rect 12 181 652 185
rect 12 161 652 165
rect 12 141 652 145
rect 12 121 652 125
rect 24 101 652 105
<< ndiffusion >>
rect -7 72 273 76
rect -7 71 277 72
rect 296 72 576 76
rect 292 71 576 72
rect -7 66 277 67
rect -7 62 76 66
rect 80 62 277 66
rect 292 66 576 67
rect 292 62 543 66
rect 547 62 576 66
rect -7 52 273 56
rect -7 51 277 52
rect 296 52 576 56
rect 292 51 576 52
rect -7 46 277 47
rect -7 42 76 46
rect 80 42 277 46
rect 292 46 576 47
rect 292 42 528 46
rect 532 42 576 46
rect 29 32 305 36
rect 29 31 309 32
rect 29 26 309 27
rect 33 22 309 26
rect -3 12 561 16
rect -7 11 561 12
rect -7 6 561 7
rect -7 2 76 6
rect 80 2 561 6
rect -3 -8 561 -4
rect -7 -9 561 -8
rect -7 -14 561 -13
rect -7 -18 312 -14
rect 316 -18 557 -14
<< pdiffusion >>
rect 12 186 648 190
rect 12 185 652 186
rect 12 180 652 181
rect 12 176 564 180
rect 568 176 652 180
rect 12 166 648 170
rect 12 165 652 166
rect 12 160 652 161
rect 12 156 554 160
rect 558 156 652 160
rect 12 146 564 150
rect 568 146 652 150
rect 12 145 652 146
rect 12 140 652 141
rect 12 136 22 140
rect 26 136 543 140
rect 547 136 652 140
rect 12 126 554 130
rect 558 126 652 130
rect 12 125 652 126
rect 12 120 652 121
rect 12 116 17 120
rect 21 116 528 120
rect 532 116 652 120
rect 24 106 648 110
rect 24 105 652 106
rect 24 100 652 101
rect 24 96 282 100
rect 286 96 652 100
<< ndcontact >>
rect 273 72 277 76
rect 292 72 296 76
rect 76 62 80 66
rect 543 62 547 66
rect 273 52 277 56
rect 292 52 296 56
rect 76 42 80 46
rect 528 42 532 46
rect 305 32 309 36
rect 29 22 33 26
rect -7 12 -3 16
rect 76 2 80 6
rect -7 -8 -3 -4
rect 312 -18 316 -14
rect 557 -18 561 -14
<< pdcontact >>
rect 648 186 652 190
rect 564 176 568 180
rect 648 166 652 170
rect 554 156 558 160
rect 564 146 568 150
rect 22 136 26 140
rect 543 136 547 140
rect 554 126 558 130
rect 17 116 21 120
rect 528 116 532 120
rect 648 106 652 110
rect 282 96 286 100
<< psubstratepcontact >>
rect -26 212 -22 216
rect -16 212 -12 216
rect -6 212 -2 216
rect 4 212 8 216
rect 14 212 18 216
rect 24 212 28 216
rect 34 212 38 216
rect 44 212 48 216
rect 54 212 58 216
rect 64 212 68 216
rect 74 212 78 216
rect 84 212 88 216
rect 94 212 98 216
rect 104 212 108 216
rect 114 212 118 216
rect 124 212 128 216
rect 134 212 138 216
rect 144 212 148 216
rect 154 212 158 216
rect 164 212 168 216
rect 174 212 178 216
rect 184 212 188 216
rect 194 212 198 216
rect 204 212 208 216
rect 214 212 218 216
rect 224 212 228 216
rect 234 212 238 216
rect 244 212 248 216
rect 254 212 258 216
rect 264 212 268 216
rect 274 212 278 216
rect 284 212 288 216
rect 294 212 298 216
rect 304 212 308 216
rect 314 212 318 216
rect 324 212 328 216
rect 334 212 338 216
rect 344 212 348 216
rect 354 212 358 216
rect 364 212 368 216
rect 374 212 378 216
rect 384 212 388 216
rect 394 212 398 216
rect 404 212 408 216
rect 414 212 418 216
rect 424 212 428 216
rect 434 212 438 216
rect 444 212 448 216
rect 454 212 458 216
rect 464 212 468 216
rect 474 212 478 216
rect 484 212 488 216
rect 494 212 498 216
rect 504 212 508 216
rect 514 212 518 216
rect 524 212 528 216
rect 534 212 538 216
rect 544 212 548 216
rect 554 212 558 216
rect 564 212 568 216
rect 574 212 578 216
rect 584 212 588 216
rect 594 212 598 216
rect 604 212 608 216
rect 614 212 618 216
rect 624 212 628 216
rect 634 212 638 216
rect 644 212 648 216
rect 654 212 658 216
rect 664 212 668 216
rect 674 212 678 216
rect 684 212 690 216
rect -26 202 -22 206
rect -7 202 -3 206
rect 686 202 690 206
rect -26 192 -22 196
rect -7 192 -3 196
rect 686 192 690 196
rect -26 182 -22 186
rect -7 182 -3 186
rect 686 182 690 186
rect -26 172 -22 176
rect -7 172 -3 176
rect 686 172 690 176
rect -26 162 -22 166
rect -7 162 -3 166
rect 686 162 690 166
rect -26 152 -22 156
rect -7 152 -3 156
rect 686 152 690 156
rect -26 142 -22 146
rect -7 142 -3 146
rect 686 142 690 146
rect -26 132 -22 136
rect -7 132 -3 136
rect 686 132 690 136
rect -26 122 -22 126
rect -7 122 -3 126
rect 686 122 690 126
rect -26 112 -22 116
rect -7 112 -3 116
rect 686 112 690 116
rect -26 102 -22 106
rect -7 102 -3 106
rect 686 102 690 106
rect -26 92 -22 96
rect -7 92 -3 96
rect 686 92 690 96
rect -26 82 -22 86
rect 686 82 690 86
rect -26 72 -22 76
rect 595 72 599 76
rect 614 72 618 76
rect 633 72 637 76
rect 652 72 656 76
rect 669 72 673 76
rect 686 72 690 76
rect -26 62 -22 66
rect 595 62 599 66
rect 614 62 618 66
rect 633 62 637 66
rect 652 62 656 66
rect 669 62 673 66
rect 686 62 690 66
rect -26 52 -22 56
rect 595 52 599 56
rect 614 52 618 56
rect 633 52 637 56
rect 652 52 656 56
rect 669 52 673 56
rect 686 52 690 56
rect -26 42 -22 46
rect 595 42 599 46
rect 614 42 618 46
rect 633 42 637 46
rect 652 42 656 46
rect 669 42 673 46
rect 686 42 690 46
rect -26 32 -22 36
rect 595 32 599 36
rect 614 32 618 36
rect 633 32 637 36
rect 652 32 656 36
rect 669 32 673 36
rect 686 32 690 36
rect -14 26 -10 30
rect -4 26 0 30
rect 6 26 10 30
rect 344 27 348 31
rect 354 27 358 31
rect 364 27 368 31
rect 374 27 378 31
rect 384 27 388 31
rect 394 27 398 31
rect 404 27 408 31
rect 414 27 418 31
rect 424 27 428 31
rect 434 27 438 31
rect 444 27 448 31
rect 454 27 458 31
rect 464 27 468 31
rect 474 27 478 31
rect 484 27 488 31
rect 494 27 498 31
rect 504 27 508 31
rect 514 27 518 31
rect 524 27 528 31
rect 534 27 538 31
rect 544 27 548 31
rect 554 27 558 31
rect 564 27 568 31
rect 574 27 578 31
rect 584 27 588 31
rect -26 22 -22 26
rect 595 22 599 26
rect 614 22 618 26
rect 633 22 637 26
rect 652 22 656 26
rect 669 22 673 26
rect 686 22 690 26
rect -26 12 -22 16
rect 595 12 599 16
rect 614 12 618 16
rect 633 12 637 16
rect 652 12 656 16
rect 669 12 673 16
rect 686 12 690 16
rect -26 2 -22 6
rect 595 2 599 6
rect 614 2 618 6
rect 633 2 637 6
rect 652 2 656 6
rect 669 2 673 6
rect 686 2 690 6
rect -26 -8 -22 -4
rect 595 -8 599 -4
rect 614 -8 618 -4
rect 633 -8 637 -4
rect 652 -8 656 -4
rect 669 -8 673 -4
rect 686 -8 690 -4
rect -26 -18 -22 -14
rect 595 -18 599 -14
rect 614 -18 618 -14
rect 633 -18 637 -14
rect 652 -18 656 -14
rect 669 -18 673 -14
rect 686 -18 690 -14
rect -26 -28 -22 -24
rect 595 -28 599 -24
rect 614 -28 618 -24
rect 633 -28 637 -24
rect 652 -28 656 -24
rect 669 -28 673 -24
rect 686 -28 690 -24
rect -26 -38 -22 -34
rect -16 -38 -12 -34
rect -6 -38 -2 -34
rect 4 -38 8 -34
rect 14 -38 18 -34
rect 24 -38 28 -34
rect 34 -38 38 -34
rect 44 -38 48 -34
rect 54 -38 58 -34
rect 64 -38 68 -34
rect 74 -38 78 -34
rect 84 -38 88 -34
rect 94 -38 98 -34
rect 104 -38 108 -34
rect 114 -38 118 -34
rect 124 -38 128 -34
rect 134 -38 138 -34
rect 144 -38 148 -34
rect 154 -38 158 -34
rect 164 -38 168 -34
rect 174 -38 178 -34
rect 184 -38 188 -34
rect 194 -38 198 -34
rect 204 -38 208 -34
rect 214 -38 218 -34
rect 224 -38 228 -34
rect 234 -38 238 -34
rect 244 -38 248 -34
rect 254 -38 258 -34
rect 264 -38 268 -34
rect 274 -38 278 -34
rect 284 -38 288 -34
rect 294 -38 298 -34
rect 304 -38 308 -34
rect 314 -38 318 -34
rect 324 -38 328 -34
rect 334 -38 338 -34
rect 344 -38 348 -34
rect 354 -38 358 -34
rect 364 -38 368 -34
rect 374 -38 378 -34
rect 384 -38 388 -34
rect 394 -38 398 -34
rect 404 -38 408 -34
rect 414 -38 418 -34
rect 424 -38 428 -34
rect 434 -38 438 -34
rect 444 -38 448 -34
rect 454 -38 458 -34
rect 464 -38 468 -34
rect 474 -38 478 -34
rect 484 -38 488 -34
rect 494 -38 498 -34
rect 504 -38 508 -34
rect 514 -38 518 -34
rect 524 -38 528 -34
rect 534 -38 538 -34
rect 544 -38 548 -34
rect 554 -38 558 -34
rect 564 -38 568 -34
rect 574 -38 578 -34
rect 584 -38 588 -34
rect 594 -38 598 -34
rect 604 -38 608 -34
rect 614 -38 618 -34
rect 628 -38 632 -34
rect 638 -38 642 -34
rect 648 -38 652 -34
rect 662 -38 666 -34
rect 672 -38 676 -34
rect 682 -38 690 -34
<< nsubstratencontact >>
rect 662 186 666 190
rect 662 176 666 180
rect 662 166 666 170
rect 662 156 666 160
rect 662 146 666 150
rect 662 136 666 140
rect 662 126 666 130
rect 662 116 666 120
rect 662 106 666 110
rect 662 96 666 100
<< polysilicon >>
rect 10 181 12 185
rect 652 181 655 185
rect 10 161 12 165
rect 652 161 655 165
rect 10 141 12 145
rect 652 141 655 145
rect 10 121 12 125
rect 652 121 655 125
rect 21 101 24 105
rect 652 101 655 105
rect -10 67 -7 71
rect 277 67 280 71
rect 289 67 292 71
rect 576 67 579 71
rect -10 47 -7 51
rect 277 47 280 51
rect 289 47 292 51
rect 576 47 579 51
rect 26 27 29 31
rect 309 27 312 31
rect -10 7 -7 11
rect 561 7 564 11
rect -10 -13 -7 -9
rect 561 -13 564 -9
<< polycontact >>
rect 6 181 10 185
rect 6 161 10 165
rect 6 141 10 145
rect 6 121 10 125
rect 17 101 21 105
rect -14 67 -10 71
rect 579 67 583 71
rect -14 47 -10 51
rect 579 47 583 51
rect 312 27 316 31
rect 564 7 568 11
rect 564 -13 568 -9
<< metal1 >>
rect -30 216 694 220
rect -30 212 -26 216
rect -22 212 -16 216
rect -12 212 -6 216
rect -2 212 4 216
rect 8 212 14 216
rect 18 212 24 216
rect 28 212 34 216
rect 38 212 44 216
rect 48 212 54 216
rect 58 212 64 216
rect 68 212 74 216
rect 78 212 84 216
rect 88 212 94 216
rect 98 212 104 216
rect 108 212 114 216
rect 118 212 124 216
rect 128 212 134 216
rect 138 212 144 216
rect 148 212 154 216
rect 158 212 164 216
rect 168 212 174 216
rect 178 212 184 216
rect 188 212 194 216
rect 198 212 204 216
rect 208 212 214 216
rect 218 212 224 216
rect 228 212 234 216
rect 238 212 244 216
rect 248 212 254 216
rect 258 212 264 216
rect 268 212 274 216
rect 278 212 284 216
rect 288 212 294 216
rect 298 212 304 216
rect 308 212 314 216
rect 318 212 324 216
rect 328 212 334 216
rect 338 212 344 216
rect 348 212 354 216
rect 358 212 364 216
rect 368 212 374 216
rect 378 212 384 216
rect 388 212 394 216
rect 398 212 404 216
rect 408 212 414 216
rect 418 212 424 216
rect 428 212 434 216
rect 438 212 444 216
rect 448 212 454 216
rect 458 212 464 216
rect 468 212 474 216
rect 478 212 484 216
rect 488 212 494 216
rect 498 212 504 216
rect 508 212 514 216
rect 518 212 524 216
rect 528 212 534 216
rect 538 212 544 216
rect 548 212 554 216
rect 558 212 564 216
rect 568 212 574 216
rect 578 212 584 216
rect 588 212 594 216
rect 598 212 604 216
rect 608 212 614 216
rect 618 212 624 216
rect 628 212 634 216
rect 638 212 644 216
rect 648 212 654 216
rect 658 212 664 216
rect 668 212 674 216
rect 678 212 684 216
rect 690 212 694 216
rect -30 208 694 212
rect -30 206 -18 208
rect -30 202 -26 206
rect -22 202 -18 206
rect -30 196 -18 202
rect -30 192 -26 196
rect -22 192 -18 196
rect -30 186 -18 192
rect -30 182 -26 186
rect -22 182 -18 186
rect -30 176 -18 182
rect -30 172 -26 176
rect -22 172 -18 176
rect -30 166 -18 172
rect -30 162 -26 166
rect -22 162 -18 166
rect -30 156 -18 162
rect -30 152 -26 156
rect -22 152 -18 156
rect -30 146 -18 152
rect -30 142 -26 146
rect -22 142 -18 146
rect -30 136 -18 142
rect -30 132 -26 136
rect -22 132 -18 136
rect -30 126 -18 132
rect -30 122 -26 126
rect -22 122 -18 126
rect -30 116 -18 122
rect -30 112 -26 116
rect -22 112 -18 116
rect -30 106 -18 112
rect -30 102 -26 106
rect -22 102 -18 106
rect -30 96 -18 102
rect -30 92 -26 96
rect -22 92 -18 96
rect -30 86 -18 92
rect -10 206 0 208
rect -10 202 -7 206
rect -3 202 0 206
rect -10 196 0 202
rect 682 206 694 208
rect 682 202 686 206
rect 690 202 694 206
rect 682 196 694 202
rect -10 192 -7 196
rect -3 192 0 196
rect -10 186 0 192
rect 658 190 670 196
rect 652 186 662 190
rect 666 186 670 190
rect -10 182 -7 186
rect -3 182 0 186
rect -10 176 0 182
rect -10 172 -7 176
rect -3 172 0 176
rect -10 166 0 172
rect -10 162 -7 166
rect -3 162 0 166
rect -10 156 0 162
rect 6 165 10 181
rect 658 180 670 186
rect 10 161 26 165
rect -10 152 -7 156
rect -3 152 0 156
rect -10 146 0 152
rect -10 142 -7 146
rect -3 142 0 146
rect -10 136 0 142
rect -10 132 -7 136
rect -3 132 0 136
rect -10 126 0 132
rect -10 122 -7 126
rect -3 122 0 126
rect -10 116 0 122
rect 6 125 10 141
rect 22 140 26 161
rect -10 112 -7 116
rect -3 112 0 116
rect -10 106 0 112
rect -10 102 -7 106
rect -3 102 0 106
rect -10 96 0 102
rect 17 105 21 116
rect -10 92 -7 96
rect -3 92 0 96
rect -10 87 0 92
rect 282 88 286 96
rect -30 82 -26 86
rect -22 82 -18 86
rect -30 76 -18 82
rect -30 72 -26 76
rect -22 72 -18 76
rect -30 66 -18 72
rect -14 71 -10 75
rect 277 72 292 76
rect -30 62 -26 66
rect -22 62 -18 66
rect -30 56 -18 62
rect -30 52 -26 56
rect -22 52 -18 56
rect -30 46 -18 52
rect -14 51 -10 55
rect -30 42 -26 46
rect -22 42 -18 46
rect -30 36 -18 42
rect -30 32 -26 36
rect -22 34 -18 36
rect 76 46 80 62
rect 277 52 292 56
rect 528 46 532 116
rect 543 66 547 136
rect 554 130 558 156
rect 564 150 568 176
rect 658 176 662 180
rect 666 176 670 180
rect 658 170 670 176
rect 652 166 662 170
rect 666 166 670 170
rect 658 160 670 166
rect 658 156 662 160
rect 666 156 670 160
rect 658 150 670 156
rect 658 146 662 150
rect 666 146 670 150
rect 658 140 670 146
rect 658 136 662 140
rect 666 136 670 140
rect 658 130 670 136
rect 658 126 662 130
rect 666 126 670 130
rect 658 120 670 126
rect 658 116 662 120
rect 666 116 670 120
rect 658 110 670 116
rect 652 106 662 110
rect 666 106 670 110
rect 658 100 670 106
rect 658 96 662 100
rect 666 96 670 100
rect 658 90 670 96
rect 682 192 686 196
rect 690 192 694 196
rect 682 186 694 192
rect 682 182 686 186
rect 690 182 694 186
rect 682 176 694 182
rect 682 172 686 176
rect 690 172 694 176
rect 682 166 694 172
rect 682 162 686 166
rect 690 162 694 166
rect 682 156 694 162
rect 682 152 686 156
rect 690 152 694 156
rect 682 146 694 152
rect 682 142 686 146
rect 690 142 694 146
rect 682 136 694 142
rect 682 132 686 136
rect 690 132 694 136
rect 682 126 694 132
rect 682 122 686 126
rect 690 122 694 126
rect 682 116 694 122
rect 682 112 686 116
rect 690 112 694 116
rect 682 106 694 112
rect 682 102 686 106
rect 690 102 694 106
rect 682 96 694 102
rect 682 92 686 96
rect 690 92 694 96
rect 682 86 694 92
rect 682 82 686 86
rect 690 82 694 86
rect 591 76 603 82
rect 591 72 595 76
rect 599 72 603 76
rect 579 51 583 67
rect 591 66 603 72
rect 591 62 595 66
rect 599 62 603 66
rect 591 56 603 62
rect 591 52 595 56
rect 599 52 603 56
rect 591 46 603 52
rect 591 42 595 46
rect 599 42 603 46
rect -22 32 16 34
rect -30 30 16 32
rect -30 26 -14 30
rect -10 26 -4 30
rect 0 26 6 30
rect 10 26 16 30
rect -30 22 -26 26
rect -22 22 16 26
rect -30 16 -18 22
rect 29 16 33 22
rect -30 12 -26 16
rect -22 12 -7 16
rect -3 12 33 16
rect -30 6 -18 12
rect -30 2 -26 6
rect -22 2 -18 6
rect 76 6 80 42
rect 305 36 315 40
rect 320 36 324 40
rect 591 36 603 42
rect 591 35 595 36
rect 338 32 595 35
rect 599 32 603 36
rect 338 31 603 32
rect -30 -4 -18 2
rect -30 -8 -26 -4
rect -22 -8 -7 -4
rect -30 -14 -18 -8
rect -30 -18 -26 -14
rect -22 -18 -18 -14
rect 312 -14 316 27
rect 338 27 344 31
rect 348 27 354 31
rect 358 27 364 31
rect 368 27 374 31
rect 378 27 384 31
rect 388 27 394 31
rect 398 27 404 31
rect 408 27 414 31
rect 418 27 424 31
rect 428 27 434 31
rect 438 27 444 31
rect 448 27 454 31
rect 458 27 464 31
rect 468 27 474 31
rect 478 27 484 31
rect 488 27 494 31
rect 498 27 504 31
rect 508 27 514 31
rect 518 27 524 31
rect 528 27 534 31
rect 538 27 544 31
rect 548 27 554 31
rect 558 27 564 31
rect 568 27 574 31
rect 578 27 584 31
rect 588 27 603 31
rect 338 26 603 27
rect 338 23 595 26
rect 591 22 595 23
rect 599 22 603 26
rect 591 16 603 22
rect 591 12 595 16
rect 599 12 603 16
rect 564 -9 568 7
rect 564 -14 568 -13
rect 561 -18 568 -14
rect 591 6 603 12
rect 591 2 595 6
rect 599 2 603 6
rect 591 -4 603 2
rect 591 -8 595 -4
rect 599 -8 603 -4
rect 591 -14 603 -8
rect 591 -18 595 -14
rect 599 -18 603 -14
rect -30 -24 -18 -18
rect -30 -28 -26 -24
rect -22 -28 -18 -24
rect -30 -30 -18 -28
rect 591 -24 603 -18
rect 591 -28 595 -24
rect 599 -28 603 -24
rect 591 -30 603 -28
rect 610 76 622 82
rect 610 72 614 76
rect 618 72 622 76
rect 610 66 622 72
rect 610 62 614 66
rect 618 62 622 66
rect 610 56 622 62
rect 610 52 614 56
rect 618 52 622 56
rect 610 46 622 52
rect 610 42 614 46
rect 618 42 622 46
rect 610 36 622 42
rect 610 32 614 36
rect 618 32 622 36
rect 610 26 622 32
rect 610 22 614 26
rect 618 22 622 26
rect 610 16 622 22
rect 610 12 614 16
rect 618 12 622 16
rect 610 6 622 12
rect 610 2 614 6
rect 618 2 622 6
rect 610 -4 622 2
rect 610 -8 614 -4
rect 618 -8 622 -4
rect 610 -14 622 -8
rect 610 -18 614 -14
rect 618 -18 622 -14
rect 610 -24 622 -18
rect 610 -28 614 -24
rect 618 -28 622 -24
rect 610 -30 622 -28
rect 629 76 641 82
rect 629 72 633 76
rect 637 72 641 76
rect 629 66 641 72
rect 629 62 633 66
rect 637 62 641 66
rect 629 56 641 62
rect 629 52 633 56
rect 637 52 641 56
rect 629 46 641 52
rect 629 42 633 46
rect 637 42 641 46
rect 629 36 641 42
rect 629 32 633 36
rect 637 32 641 36
rect 629 26 641 32
rect 629 22 633 26
rect 637 22 641 26
rect 629 16 641 22
rect 629 12 633 16
rect 637 12 641 16
rect 629 6 641 12
rect 629 2 633 6
rect 637 2 641 6
rect 629 -4 641 2
rect 629 -8 633 -4
rect 637 -8 641 -4
rect 629 -14 641 -8
rect 629 -18 633 -14
rect 637 -18 641 -14
rect 629 -24 641 -18
rect 629 -28 633 -24
rect 637 -28 641 -24
rect 629 -30 641 -28
rect 648 76 660 82
rect 648 72 652 76
rect 656 72 660 76
rect 648 66 660 72
rect 648 62 652 66
rect 656 62 660 66
rect 648 56 660 62
rect 648 52 652 56
rect 656 52 660 56
rect 648 46 660 52
rect 648 42 652 46
rect 656 42 660 46
rect 648 36 660 42
rect 648 32 652 36
rect 656 32 660 36
rect 648 26 660 32
rect 648 22 652 26
rect 656 22 660 26
rect 648 16 660 22
rect 648 12 652 16
rect 656 12 660 16
rect 648 6 660 12
rect 648 2 652 6
rect 656 2 660 6
rect 648 -4 660 2
rect 648 -8 652 -4
rect 656 -8 660 -4
rect 648 -14 660 -8
rect 648 -18 652 -14
rect 656 -18 660 -14
rect 648 -24 660 -18
rect 648 -28 652 -24
rect 656 -28 660 -24
rect 648 -30 660 -28
rect 665 76 677 82
rect 665 72 669 76
rect 673 72 677 76
rect 665 66 677 72
rect 665 62 669 66
rect 673 62 677 66
rect 665 56 677 62
rect 665 52 669 56
rect 673 52 677 56
rect 665 46 677 52
rect 665 42 669 46
rect 673 42 677 46
rect 665 36 677 42
rect 665 32 669 36
rect 673 32 677 36
rect 665 26 677 32
rect 665 22 669 26
rect 673 22 677 26
rect 665 16 677 22
rect 665 12 669 16
rect 673 12 677 16
rect 665 6 677 12
rect 665 2 669 6
rect 673 2 677 6
rect 665 -4 677 2
rect 665 -8 669 -4
rect 673 -8 677 -4
rect 665 -14 677 -8
rect 665 -18 669 -14
rect 673 -18 677 -14
rect 665 -24 677 -18
rect 665 -28 669 -24
rect 673 -28 677 -24
rect 665 -30 677 -28
rect 682 76 694 82
rect 682 72 686 76
rect 690 72 694 76
rect 682 66 694 72
rect 682 62 686 66
rect 690 62 694 66
rect 682 56 694 62
rect 682 52 686 56
rect 690 52 694 56
rect 682 46 694 52
rect 682 42 686 46
rect 690 42 694 46
rect 682 36 694 42
rect 682 32 686 36
rect 690 32 694 36
rect 682 26 694 32
rect 682 22 686 26
rect 690 22 694 26
rect 682 16 694 22
rect 682 12 686 16
rect 690 12 694 16
rect 682 6 694 12
rect 682 2 686 6
rect 690 2 694 6
rect 682 -4 694 2
rect 682 -8 686 -4
rect 690 -8 694 -4
rect 682 -14 694 -8
rect 682 -18 686 -14
rect 690 -18 694 -14
rect 682 -24 694 -18
rect 682 -28 686 -24
rect 690 -28 694 -24
rect 682 -30 694 -28
rect -30 -34 694 -30
rect -30 -38 -26 -34
rect -22 -38 -16 -34
rect -12 -38 -6 -34
rect -2 -38 4 -34
rect 8 -38 14 -34
rect 18 -38 24 -34
rect 28 -38 34 -34
rect 38 -38 44 -34
rect 48 -38 54 -34
rect 58 -38 64 -34
rect 68 -38 74 -34
rect 78 -38 84 -34
rect 88 -38 94 -34
rect 98 -38 104 -34
rect 108 -38 114 -34
rect 118 -38 124 -34
rect 128 -38 134 -34
rect 138 -38 144 -34
rect 148 -38 154 -34
rect 158 -38 164 -34
rect 168 -38 174 -34
rect 178 -38 184 -34
rect 188 -38 194 -34
rect 198 -38 204 -34
rect 208 -38 214 -34
rect 218 -38 224 -34
rect 228 -38 234 -34
rect 238 -38 244 -34
rect 248 -38 254 -34
rect 258 -38 264 -34
rect 268 -38 274 -34
rect 278 -38 284 -34
rect 288 -38 294 -34
rect 298 -38 304 -34
rect 308 -38 314 -34
rect 318 -38 324 -34
rect 328 -38 334 -34
rect 338 -38 344 -34
rect 348 -38 354 -34
rect 358 -38 364 -34
rect 368 -38 374 -34
rect 378 -38 384 -34
rect 388 -38 394 -34
rect 398 -38 404 -34
rect 408 -38 414 -34
rect 418 -38 424 -34
rect 428 -38 434 -34
rect 438 -38 444 -34
rect 448 -38 454 -34
rect 458 -38 464 -34
rect 468 -38 474 -34
rect 478 -38 484 -34
rect 488 -38 494 -34
rect 498 -38 504 -34
rect 508 -38 514 -34
rect 518 -38 524 -34
rect 528 -38 534 -34
rect 538 -38 544 -34
rect 548 -38 554 -34
rect 558 -38 564 -34
rect 568 -38 574 -34
rect 578 -38 584 -34
rect 588 -38 594 -34
rect 598 -38 604 -34
rect 608 -38 614 -34
rect 618 -38 628 -34
rect 632 -38 638 -34
rect 642 -38 648 -34
rect 652 -38 662 -34
rect 666 -38 672 -34
rect 676 -38 682 -34
rect 690 -38 694 -34
rect -30 -42 694 -38
<< m2contact >>
rect 281 83 286 88
rect 315 36 320 41
<< metal2 >>
rect 282 41 286 83
rect 282 37 315 41
<< labels >>
rlabel metal1 7 134 7 134 3 b2
rlabel metal1 530 86 530 86 3 d4
rlabel metal1 545 86 545 86 3 d3
rlabel metal1 566 154 566 154 3 d5
rlabel metal1 556 133 556 133 3 d6
rlabel metal1 580 59 580 59 3 b1
rlabel metal1 566 0 566 0 3 ref
rlabel metal1 322 38 322 38 3 out
rlabel metal1 -12 53 -12 53 3 inp
rlabel metal1 -12 73 -12 73 3 inn
rlabel metal1 78 39 78 39 3 d9
rlabel metal1 278 74 278 74 3 d1
rlabel metal1 279 54 279 54 3 d2
rlabel metal1 -13 -6 -13 -6 3 gnd!
rlabel metal1 655 108 655 108 3 vdd!
<< end >>
