* SPICE3 file created from telescopic.ext - technology: scmos

.option scale=0.09u

M1000 d4 b1 d2 gnd CMOSN w=284 l=4
+  ad=1420 pd=578 as=2840 ps=1156
M1001 d4 b2 d6 vdd CMOSP w=568 l=4
+  ad=2840 pd=1146 as=5680 ps=2292
M1002 gnd ref out gnd CMOSN w=316 l=4
+  ad=7260 pd=2934 as=1580 ps=642
M1003 d6 d3 vdd vdd CMOSP w=568 l=4
+  ad=0 pd=0 as=8460 ps=3414
M1004 d3 b1 d1 gnd CMOSN w=284 l=4
+  ad=1420 pd=578 as=2840 ps=1156
M1005 d9 inp d2 gnd CMOSN w=284 l=4
+  ad=5680 pd=2302 as=0 ps=0
M1006 ref ref gnd gnd CMOSN w=568 l=4
+  ad=2840 pd=1146 as=0 ps=0
M1007 d3 b2 d5 vdd CMOSP w=568 l=4
+  ad=2840 pd=1146 as=5680 ps=2292
M1008 d9 inn d1 gnd CMOSN w=284 l=4
+  ad=0 pd=0 as=0 ps=0
M1009 d5 d3 vdd vdd CMOSP w=568 l=4
+  ad=0 pd=0 as=0 ps=0
M1010 out d4 vdd vdd CMOSP w=556 l=4
+  ad=2780 pd=1122 as=0 ps=0
M1011 d9 ref gnd gnd CMOSN w=568 l=4
+  ad=0 pd=0 as=0 ps=0
C0 d6 vdd 0.04fF
C1 gnd ref 0.04fF
C2 d5 d3 0.12fF
C3 d4 d1 0.02fF
C4 d5 vdd 0.06fF
C5 d4 gnd 0.02fF
C6 d4 d3 0.14fF
C7 d4 vdd 0.21fF
C8 b2 gnd 0.16fF
C9 b2 d3 0.21fF
C10 d3 d1 0.02fF
C11 out d9 0.02fF
C12 d9 inp 0.10fF
C13 b2 vdd 0.23fF
C14 d3 gnd 0.16fF
C15 d3 vdd 0.35fF
C16 d9 ref 0.23fF
C17 b1 d4 0.21fF
C18 out ref 0.03fF
C19 d9 d2 0.02fF
C20 out d4 0.02fF
C21 d6 d5 0.13fF
C22 out d2 0.09fF
C23 gnd d9 0.04fF
C24 b1 d3 0.10fF
C25 out d1 0.11fF
C26 gnd inp 0.08fF
C27 out d3 0.02fF
C28 d6 b2 0.10fF
C29 out vdd 0.02fF
C30 gnd inn 0.08fF
C31 d6 d3 0.15fF
C32 d4 d2 0.02fF
C33 d9 gnd 0.06fF
C34 inp gnd 0.13fF
C35 inn gnd 0.13fF
C36 ref gnd 0.49fF
C37 d2 gnd 0.06fF
C38 d1 gnd 0.06fF
C39 b1 gnd 0.04fF
C40 out gnd 0.91fF
C41 d6 gnd 0.00fF
C42 d5 gnd 0.00fF
C43 d4 gnd 0.07fF
C44 b2 gnd 0.04fF
C45 d3 gnd 0.09fF
C46 gnd gnd 12.02fF
C47 vdd gnd 63.16fF
