* Telescopic
.include TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param length=0.36u

.param width_1234={0.36*71u}
.param width_5678={0.36*160u}
.param width_910={0.36*142u}
.param width_11={0.36*157u}
.param width_12={0.36*70u}

.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
Iref gnd ref 400u
Vb1 b1 gnd 1.4
Vb2 b2 gnd 0.75

*op
*vinp inp gnd 0.9

* Transient and AC
* vinp inp gnd dc 0.9 ac 0.01m sin(0.9 0.01m 10k 0 0 0)

* Slew Rate
*vinp inp gnd pulse(1 0 -1n 100p 100p 500n 1u)

* Offset
vinp inp gnd 0.9

*vinp inp gnd dc 0.9 ac 0.6 sin(0.9 0.6 10k 0 0 0)

Cc k inn 2p
Rs d4 k 1k

M1      d1     inn      d9     gnd  CMOSN   W={width_1234}   L={length}
+ AS={5*width_1234*LAMBDA} PS={10*LAMBDA+2*width_1234} AD={5*width_1234*LAMBDA} PD={10*LAMBDA+2*width_1234}
M2      d2     inp      d9     gnd  CMOSN   W={width_1234}   L={length}
+ AS={5*width_1234*LAMBDA} PS={10*LAMBDA+2*width_1234} AD={5*width_1234*LAMBDA} PD={10*LAMBDA+2*width_1234}
M3      d3     b1       d1    gnd  CMOSN   W={width_1234}   L={length}
+ AS={5*width_1234*LAMBDA} PS={10*LAMBDA+2*width_1234} AD={5*width_1234*LAMBDA} PD={10*LAMBDA+2*width_1234}
M4      d4     b1       d2    gnd  CMOSN   W={width_1234}   L={length}
+ AS={5*width_1234*LAMBDA} PS={10*LAMBDA+2*width_1234} AD={5*width_1234*LAMBDA} PD={10*LAMBDA+2*width_1234}
M5      d3     b2      d5     vdd  CMOSP   W={width_5678}   L={length}
+ AS={5*width_5678*LAMBDA} PS={10*LAMBDA+2*width_5678} AD={5*width_5678*LAMBDA} PD={10*LAMBDA+2*width_5678}
M6      d4     b2      d6     vdd  CMOSP   W={width_5678}   L={length}
+ AS={5*width_5678*LAMBDA} PS={10*LAMBDA+2*width_5678} AD={5*width_5678*LAMBDA} PD={10*LAMBDA+2*width_5678}
M7      d5     d3       vdd    vdd  CMOSP   W={width_5678}   L={length}
+ AS={5*width_5678*LAMBDA} PS={10*LAMBDA+2*width_5678} AD={5*width_5678*LAMBDA} PD={10*LAMBDA+2*width_5678}
M8      d6     d3       vdd    vdd  CMOSP   W={width_5678}   L={length}
+ AS={5*width_5678*LAMBDA} PS={10*LAMBDA+2*width_5678} AD={5*width_5678*LAMBDA} PD={10*LAMBDA+2*width_5678}


M9      d9    ref      gnd    gnd  CMOSN   W={width_910}   L={length}
+ AS={5*width_910*LAMBDA} PS={10*LAMBDA+2*width_910} AD={5*width_910*LAMBDA} PD={10*LAMBDA+2*width_910}
M10      ref     ref     gnd     gnd  CMOSN   W={width_910}   L={length}
+ AS={5*width_910*LAMBDA} PS={10*LAMBDA+2*width_910} AD={5*width_910*LAMBDA} PD={10*LAMBDA+2*width_910}

M11      inn    d4       vdd    vdd  CMOSP   W={width_11}   L={length}
+ AS={5*width_11*LAMBDA} PS={10*LAMBDA+2*width_11} AD={5*width_11*LAMBDA} PD={10*LAMBDA+2*width_11}
M12      inn    ref      gnd     gnd  CMOSN   W={width_12}   L={length}
+ AS={5*width_12*LAMBDA} PS={10*LAMBDA+2*width_12} AD={5*width_12*LAMBDA} PD={10*LAMBDA+2*width_12}

*.tran 1u 1m
*.op
*.ac dec 10 1 1000Meg
*.dc vinp 0 1.8 0.01


* Slew rate & Offset
*.tran 0.001u 1u

.control
run

set hcopypscolor = 1
set color0=white
set color1=black

*plot v(inn) v(inp)

*plot v(inp) v(inn) deriv(v(inn))
*plot v(inp)-v(inn)

*fourier 10k v(inp)-v(inn)
*fourier 10k v(inn)

*plot v(inn)/v(inp)
*plot 180/PI*phase(v(inn)/(v(inp)))

*plot (db(v(inn))-db(v(inp))) 
*plot 180/PI*phase(v(inn)/(v(inp)))

* Slew rate
plot v(inp) V(inn)
*plot deriv(v(inn))

* PSRR
*plot v(inn)
*plot v(inn)/v(vdd)
*plot (db(v(inn))-db(v(vdd)))

* ICMR 
*plot v(inn)
*plot deriv(v(inn))

.endc
