* SPICE3 file created from telescopic.ext - technology: scmos

.option scale=0.09u

M1000 d4 b1 d2 gnd CMOSN w=284 l=4
+  ad=1420 pd=578 as=2840 ps=1156
M1001 d4 b2 d6 vdd CMOSP w=640 l=4
+  ad=3200 pd=1290 as=6400 ps=2580
M1002 gnd ref out gnd CMOSN w=316 l=4
+  ad=7260 pd=2934 as=1580 ps=642
M1003 d6 d3 vdd vdd CMOSP w=640 l=4
+  ad=0 pd=0 as=9540 ps=3846
M1004 d3 b1 d1 gnd CMOSN w=284 l=4
+  ad=1420 pd=578 as=2840 ps=1156
M1005 d9 inp d2 gnd CMOSN w=284 l=4
+  ad=5680 pd=2302 as=0 ps=0
M1006 ref ref gnd gnd CMOSN w=568 l=4
+  ad=2840 pd=1146 as=0 ps=0
M1007 d3 b2 d5 vdd CMOSP w=640 l=4
+  ad=3200 pd=1290 as=6400 ps=2580
M1008 d9 inn d1 gnd CMOSN w=284 l=4
+  ad=0 pd=0 as=0 ps=0
M1009 d5 d3 vdd vdd CMOSP w=640 l=4
+  ad=0 pd=0 as=0 ps=0
M1010 out d4 vdd vdd CMOSP w=628 l=4
+  ad=3140 pd=1266 as=0 ps=0
M1011 d9 ref gnd gnd CMOSN w=568 l=4
+  ad=0 pd=0 as=0 ps=0
C0 out d9 0.02fF
C1 d4 out 0.02fF
C2 d5 d6 0.13fF
C3 d3 d1 0.02fF
C4 vdd d6 0.04fF
C5 d4 b1 0.21fF
C6 vdd out 0.02fF
C7 d4 d1 0.02fF
C8 d2 d9 0.02fF
C9 d4 d2 0.02fF
C10 ref d9 0.23fF
C11 d3 b2 0.21fF
C12 out d1 0.11fF
C13 d3 d4 0.14fF
C14 inp d9 0.10fF
C15 out d2 0.09fF
C16 d3 d5 0.12fF
C17 gnd ref 0.04fF
C18 vdd d3 0.35fF
C19 out ref 0.03fF
C20 d3 d6 0.15fF
C21 gnd inn 0.08fF
C22 gnd d3 0.16fF
C23 vdd b2 0.23fF
C24 gnd inp 0.08fF
C25 d3 out 0.02fF
C26 b2 d6 0.10fF
C27 vdd d4 0.21fF
C28 gnd b2 0.16fF
C29 d3 b1 0.10fF
C30 gnd d9 0.04fF
C31 vdd d5 0.06fF
C32 gnd d4 0.02fF
C33 d9 gnd 0.06fF
C34 inp gnd 0.13fF
C35 inn gnd 0.13fF
C36 ref gnd 0.49fF
C37 d2 gnd 0.06fF
C38 d1 gnd 0.06fF
C39 b1 gnd 0.04fF
C40 out gnd 0.91fF
C41 d6 gnd 0.00fF
C42 d5 gnd 0.00fF
C43 d4 gnd 0.07fF
C44 b2 gnd 0.04fF
C45 d3 gnd 0.09fF
C46 gnd gnd 15.15fF
C47 vdd gnd 70.82fF
